//`timescale 1ns / 1ps

//module full_adder(
//    input x, y, z,
//    output c, s
//    );
    
//    // s = xy' + x'y
//    assign s = (x & ~y) | (~x & y);
    
//    // c = xy
//    assign c = x & y;
//endmodule
